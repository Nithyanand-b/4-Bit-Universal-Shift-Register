module four_bit_USR (
    input wire clk,
    input wire rst,
    input wire [1:0] mode,
    input wire [3:0] data_in,
    input wire serial_in,
    output reg [3:0] data_out
);

always @(posedge clk or posedge rst) begin
    if (rst)
        data_out <= 4'b0000;
    else begin
        case (mode)
            2'b00: data_out <= data_out; // Hold
            2'b01: data_out <= {serial_in, data_out[3:1]}; // Shift right
            2'b10: data_out <= {data_out[2:0], serial_in}; // Shift left
            2'b11: data_out <= data_in; // Parallel load
        endcase
    end
end

endmodule
